library verilog;
use verilog.vl_types.all;
entity key_loader_struct_vlg_vec_tst is
end key_loader_struct_vlg_vec_tst;
