library verilog;
use verilog.vl_types.all;
entity matrix_mult_struct_vlg_vec_tst is
end matrix_mult_struct_vlg_vec_tst;
