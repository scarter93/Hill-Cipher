library verilog;
use verilog.vl_types.all;
entity key_inverter_vlg_vec_tst is
end key_inverter_vlg_vec_tst;
