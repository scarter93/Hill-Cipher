library verilog;
use verilog.vl_types.all;
entity hill_cipher_vlg_vec_tst is
end hill_cipher_vlg_vec_tst;
